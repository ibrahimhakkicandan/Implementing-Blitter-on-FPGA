module intf_axi4 (



);
